module day04

const pattern_1d = [`X`, `M`, `A`, `S`]

const pattern_1d_reverse = [`S`, `A`, `M`, `X`]

const pattern_2d = [
	[`X`, ` `, ` `, ` `],
	[` `, `M`, ` `, ` `],
	[` `, ` `, `A`, ` `],
	[` `, ` `, ` `, `S`],
]

const pattern_2d_reverse = [
	[`S`, ` `, ` `, ` `],
	[` `, `A`, ` `, ` `],
	[` `, ` `, `M`, ` `],
	[` `, ` `, ` `, `X`],
]
