module day04

const pattern_1d = [`X`, `M`, `A`, `S`]

const pattern_1d_reverse = [`S`, `A`, `M`, `X`]

const pattern_2d = [
	[`X`, ` `, ` `, ` `],
	[` `, `M`, ` `, ` `],
	[` `, ` `, `A`, ` `],
	[` `, ` `, ` `, `S`],
]

const pattern_2d_reverse = [
	[`S`, ` `, ` `, ` `],
	[` `, `A`, ` `, ` `],
	[` `, ` `, `M`, ` `],
	[` `, ` `, ` `, `X`],
]

const pattern_2_2d = [
	[`M`, ` `, `S`],
	[` `, `A`, ` `],
	[`M`, ` `, `S`],
]

const pattern_2_2d_2 = [
	[`S`, ` `, `S`],
	[` `, `A`, ` `],
	[`M`, ` `, `M`],
]

const pattern_2_2d_3 = [
	[`M`, ` `, `M`],
	[` `, `A`, ` `],
	[`S`, ` `, `S`],
]

const pattern_2_2d_4 = [
	[`S`, ` `, `M`],
	[` `, `A`, ` `],
	[`S`, ` `, `M`],
]
